module knight_attack2_50_64_IVT_example (
	input logic vga_clk,
	input logic [9:0] DrawX, DrawY,
	input logic blank,
	output logic [3:0] red, green, blue
);

logic [11:0] rom_address;
logic [2:0] rom_q;

logic [3:0] palette_red, palette_green, palette_blue;

logic negedge_vga_clk;

// read from ROM on negedge, set pixel on posedge
assign negedge_vga_clk = ~vga_clk;

// address into the rom = (x*xDim)/640 + ((y*yDim)/480) * xDim
// this will stretch out the sprite across the entire screen
assign rom_address = ((DrawX * 50) / 640) + (((DrawY * 64) / 480) * 50);

always_ff @ (posedge vga_clk) begin
	red <= 4'h0;
	green <= 4'h0;
	blue <= 4'h0;

	if (blank) begin
		red <= palette_red;
		green <= palette_green;
		blue <= palette_blue;
	end
end

knight_attack2_50_64_IVT_rom knight_attack2_50_64_IVT_rom (
	.clock   (negedge_vga_clk),
	.address (rom_address_at2I),
	.q       (rom_q_at2I)
);

knight_attack2_50_64_IVT_palette knight_attack2_50_64_IVT_palette (
	.index (rom_q_at2I),
	.red   (palette_red_at2I),
	.green (palette_green_at2I),
	.blue  (palette_blue_at2I)
);

endmodule
